Library ieee;
USE ieee.std_logic_1164.all;

package lab1_1_package IS

	component lab1_1
		PORT (w, x, y, z : IN STD_LOGIC;
				a, b, c, d, e, f, g : OUT STD_LOGIC);
	end component;
	
END lab1_1_package;



